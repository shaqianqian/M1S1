library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity SORT8 is
    Port ( U1 : in  STD_LOGIC_VECTOR (8 downto 0);
           U2 : in  STD_LOGIC_VECTOR (8 downto 0);
           U3 : in  STD_LOGIC_VECTOR (8 downto 0);
           U4 : in  STD_LOGIC_VECTOR (8 downto 0);
           U5 : in  STD_LOGIC_VECTOR (8 downto 0);
           U6 : in  STD_LOGIC_VECTOR (8 downto 0);
           U7 : in  STD_LOGIC_VECTOR (8 downto 0);
           U8 : in  STD_LOGIC_VECTOR (8 downto 0);
           Z1 : out  STD_LOGIC_VECTOR (8 downto 0);
           Z2 : out  STD_LOGIC_VECTOR (8 downto 0);
           Z3 : out  STD_LOGIC_VECTOR (8 downto 0);
           Z4 : out  STD_LOGIC_VECTOR (8 downto 0);
           Z5 : out  STD_LOGIC_VECTOR (8 downto 0);
           Z6 : out  STD_LOGIC_VECTOR (8 downto 0);
           Z7 : out  STD_LOGIC_VECTOR (8 downto 0);
           Z8 : out  STD_LOGIC_VECTOR (8 downto 0));
end SORT8;

architecture Behavioral of SORT8 is

begin


end Behavioral;

